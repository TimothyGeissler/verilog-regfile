module test1_tb();
    
endmodule